library verilog;
use verilog.vl_types.all;
entity Instruction_system_vlg_vec_tst is
end Instruction_system_vlg_vec_tst;
