library verilog;
use verilog.vl_types.all;
entity CPU_vlg_vec_tst is
end CPU_vlg_vec_tst;
